	 module hpi_io_intf( input [1:0]  from_sw_address,
								output[15:0] from_sw_data_in,
								input [15:0] from_sw_data_out,
								input		 	 from_sw_r,from_sw_w,from_sw_cs,
								inout [15:0] OTG_DATA,    
								output[1:0]	 OTG_ADDR,    
								output		 OTG_RD_N, OTG_WR_N, OTG_CS_N, OTG_RST_N, 
								input 		 OTG_INT, Clk, Reset);
								
logic [15:0] tmp_data;
logic from_sw_int; 

//Fill in the blanks below. 
// ~~~ All following ocmmented lines are commented for the sake of compilation (Jacob)
// assign OTG_RST_N = 
// assign OTG_DATA = //Should be tristated

//always_ff @ (posedge Clk or posedge Reset)
//begin
//	if(Reset)
//	begin
//		tmp_data 		<= 
//		OTG_ADDR 		<=	2b'0;
//		OTG_RD_N 		<= 0;
//		OTG_WR_N 		<= 0;
//		OTG_CS_N 		<= 0;
//		from_sw_data_in<= 0;
//		from_sw_int 	<= 
//	end
//	else 
//	begin
//		tmp_data 		<= 
//		OTG_ADDR 		<= 
//		OTG_RD_N			<= 
//		OTG_WR_N			<= 
//		OTG_CS_N			<= 
//		from_sw_data_in<= 
//		from_sw_int 	<= 
//	end
//end
endmodule 