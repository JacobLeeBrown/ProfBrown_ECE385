module  circle(output [29:0][29:0] c);
	assign c[0]  = 30'b000000000001111111100000000000;
	assign c[1]  = 30'b000000001110000000011100000000;
	assign c[2]  = 30'b000000010000000000000010000000;
	assign c[3]  = 30'b000001100000000000000001100000;
	assign c[4]  = 30'b000010000000000000000000010000;
	assign c[5]  = 30'b000100000000000000000000001000;
	assign c[6]  = 30'b000100000000000000000000001000;
	assign c[7]  = 30'b001000000000000000000000000100;
	assign c[8]  = 30'b010000000000000000000000000010;
	assign c[9]  = 30'b010000000000000000000000000010;
	assign c[10] = 30'b010000000000000000000000000010;
	assign c[11] = 30'b100000000000000000000000000001;
	assign c[12] = 30'b100000000000000000000000000001;
	assign c[13] = 30'b100000000000000000000000000001;
	assign c[14] = 30'b100000000000000000000000000001;
	assign c[15] = 30'b100000000000000000000000000001;
	assign c[16] = 30'b100000000000000000000000000001;
	assign c[17] = 30'b100000000000000000000000000001;
	assign c[18] = 30'b100000000000000000000000000001;
	assign c[19] = 30'b010000000000000000000000000010;
	assign c[20] = 30'b010000000000000000000000000010;
	assign c[21] = 30'b010000000000000000000000000010;
	assign c[22] = 30'b001000000000000000000000000100;
	assign c[23] = 30'b000100000000000000000000001000;
	assign c[24] = 30'b000100000000000000000000001000;
	assign c[25] = 30'b000010000000000000000000010000;
	assign c[26] = 30'b000001100000000000000001100000;
	assign c[27] = 30'b000000010000000000000010000000;
	assign c[28] = 30'b000000001110000000011100000000;
	assign c[29] = 30'b000000000001111111100000000000;
endmodule
