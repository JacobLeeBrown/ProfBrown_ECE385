module testbench();

timeunit 10ns;	// Half clock cycle at 50 MHz
// This is the amount of time represented by #1 
timeprecision 1ns;

// These signals are internal because the processor will be 
// instantiated as a submodule in testbench.
logic [15:0] S;
logic Clk = 0;
logic Reset, Run, Continue;
logic [11:0] LED;
logic [6:0]  HEX0, HEX1, HEX2, HEX3;
logic  CE, UB, LB, OE, WE;
logic [19:0] ADDR;
logic [15:0] Data;

// Instantiating the Processor
slc3 Big_Papa(.*);	

// Toggle the clock
// #1 means wait for a delay of 1 timeunit
always begin : CLOCK_GENERATION
#1 Clk = ~Clk;
end

initial begin: CLOCK_INITIALIZATION
    Clk = 0;
end 

// Testing begins here
// The initial block is not synthesizable
// Everything happens sequentially inside an initial block as in a software program
initial begin: TEST_VECTORS
Reset = 0;
Run = 1;
Continue = 1;

#2 Reset = 1;

// #2 ADDR = 16'hFFFF;
// #2 S = 16'b0000000001011010;	// x005A
#2 S = 16'b0000000000000011;	// x0003

#2 Run = 0;
#2 Run = 1;
/*
#6 S = 16'b1100110011001100;
#4 S = 16'b1010101010101010;
#4 S = 16'b0000111100001111;
#4 S = 16'b1111000011110000;
#4 S = 16'b0001001000110100;
*/
#10 Continue = ~Continue;
#2 Continue = ~Continue;

#10 Continue = ~Continue;
#2 Continue = ~Continue;

#10 Continue = ~Continue;
#2 Continue = ~Continue;

#10 Continue = ~Continue;
#2 Continue = ~Continue;
end
endmodule
